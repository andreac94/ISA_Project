library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity DADDA_24 is
	port (M1, M2 : in  std_logic_vector(23 downto 0);
	      PROD   : out std_logic_vector(47 downto 0)
	);
end DADDA_24;

architecture arch of DADDA_24 is

	component HA
		port (A, B : in  std_logic;
		      S, C : out std_logic
		);
	end component;

	component FA
		port (A, B, C_in : in  std_logic;
		      S, C_out   : out std_logic
		);
	end component;
	
	component ROUNDING_AND_OVF_UNIT
		generic (N : natural);
		port (I : in  std_logic_vector(2*N-1 downto 0);
		      O : out std_logic_vector(  N-1 downto 0)
		);
	end component;

	-- SIGNALS
	signal pp              : std_logic_vector(575 downto 0);
	signal sum             : std_logic_vector(505 downto 0);
	signal carry           : std_logic_vector(505 downto 0);
	signal final_adder_op1 : std_logic_vector(46 downto 0);
	signal final_adder_op2 : std_logic_vector(46 downto 0);
	signal final_adder_sum : integer;

begin
	-- PARTIAL PRODUCTS
	pp(0) <= M1(0) and M2(0);
	pp(1) <= M1(0) and M2(1);
	pp(2) <= M1(0) and M2(2);
	pp(3) <= M1(0) and M2(3);
	pp(4) <= M1(0) and M2(4);
	pp(5) <= M1(0) and M2(5);
	pp(6) <= M1(0) and M2(6);
	pp(7) <= M1(0) and M2(7);
	pp(8) <= M1(0) and M2(8);
	pp(9) <= M1(0) and M2(9);
	pp(10) <= M1(0) and M2(10);
	pp(11) <= M1(0) and M2(11);
	pp(12) <= M1(0) and M2(12);
	pp(13) <= M1(0) and M2(13);
	pp(14) <= M1(0) and M2(14);
	pp(15) <= M1(0) and M2(15);
	pp(16) <= M1(0) and M2(16);
	pp(17) <= M1(0) and M2(17);
	pp(18) <= M1(0) and M2(18);
	pp(19) <= M1(0) and M2(19);
	pp(20) <= M1(0) and M2(20);
	pp(21) <= M1(0) and M2(21);
	pp(22) <= M1(0) and M2(22);
	pp(23) <= M1(0) and M2(23);
	pp(24) <= M1(1) and M2(0);
	pp(25) <= M1(1) and M2(1);
	pp(26) <= M1(1) and M2(2);
	pp(27) <= M1(1) and M2(3);
	pp(28) <= M1(1) and M2(4);
	pp(29) <= M1(1) and M2(5);
	pp(30) <= M1(1) and M2(6);
	pp(31) <= M1(1) and M2(7);
	pp(32) <= M1(1) and M2(8);
	pp(33) <= M1(1) and M2(9);
	pp(34) <= M1(1) and M2(10);
	pp(35) <= M1(1) and M2(11);
	pp(36) <= M1(1) and M2(12);
	pp(37) <= M1(1) and M2(13);
	pp(38) <= M1(1) and M2(14);
	pp(39) <= M1(1) and M2(15);
	pp(40) <= M1(1) and M2(16);
	pp(41) <= M1(1) and M2(17);
	pp(42) <= M1(1) and M2(18);
	pp(43) <= M1(1) and M2(19);
	pp(44) <= M1(1) and M2(20);
	pp(45) <= M1(1) and M2(21);
	pp(46) <= M1(1) and M2(22);
	pp(47) <= M1(1) and M2(23);
	pp(48) <= M1(2) and M2(0);
	pp(49) <= M1(2) and M2(1);
	pp(50) <= M1(2) and M2(2);
	pp(51) <= M1(2) and M2(3);
	pp(52) <= M1(2) and M2(4);
	pp(53) <= M1(2) and M2(5);
	pp(54) <= M1(2) and M2(6);
	pp(55) <= M1(2) and M2(7);
	pp(56) <= M1(2) and M2(8);
	pp(57) <= M1(2) and M2(9);
	pp(58) <= M1(2) and M2(10);
	pp(59) <= M1(2) and M2(11);
	pp(60) <= M1(2) and M2(12);
	pp(61) <= M1(2) and M2(13);
	pp(62) <= M1(2) and M2(14);
	pp(63) <= M1(2) and M2(15);
	pp(64) <= M1(2) and M2(16);
	pp(65) <= M1(2) and M2(17);
	pp(66) <= M1(2) and M2(18);
	pp(67) <= M1(2) and M2(19);
	pp(68) <= M1(2) and M2(20);
	pp(69) <= M1(2) and M2(21);
	pp(70) <= M1(2) and M2(22);
	pp(71) <= M1(2) and M2(23);
	pp(72) <= M1(3) and M2(0);
	pp(73) <= M1(3) and M2(1);
	pp(74) <= M1(3) and M2(2);
	pp(75) <= M1(3) and M2(3);
	pp(76) <= M1(3) and M2(4);
	pp(77) <= M1(3) and M2(5);
	pp(78) <= M1(3) and M2(6);
	pp(79) <= M1(3) and M2(7);
	pp(80) <= M1(3) and M2(8);
	pp(81) <= M1(3) and M2(9);
	pp(82) <= M1(3) and M2(10);
	pp(83) <= M1(3) and M2(11);
	pp(84) <= M1(3) and M2(12);
	pp(85) <= M1(3) and M2(13);
	pp(86) <= M1(3) and M2(14);
	pp(87) <= M1(3) and M2(15);
	pp(88) <= M1(3) and M2(16);
	pp(89) <= M1(3) and M2(17);
	pp(90) <= M1(3) and M2(18);
	pp(91) <= M1(3) and M2(19);
	pp(92) <= M1(3) and M2(20);
	pp(93) <= M1(3) and M2(21);
	pp(94) <= M1(3) and M2(22);
	pp(95) <= M1(3) and M2(23);
	pp(96) <= M1(4) and M2(0);
	pp(97) <= M1(4) and M2(1);
	pp(98) <= M1(4) and M2(2);
	pp(99) <= M1(4) and M2(3);
	pp(100) <= M1(4) and M2(4);
	pp(101) <= M1(4) and M2(5);
	pp(102) <= M1(4) and M2(6);
	pp(103) <= M1(4) and M2(7);
	pp(104) <= M1(4) and M2(8);
	pp(105) <= M1(4) and M2(9);
	pp(106) <= M1(4) and M2(10);
	pp(107) <= M1(4) and M2(11);
	pp(108) <= M1(4) and M2(12);
	pp(109) <= M1(4) and M2(13);
	pp(110) <= M1(4) and M2(14);
	pp(111) <= M1(4) and M2(15);
	pp(112) <= M1(4) and M2(16);
	pp(113) <= M1(4) and M2(17);
	pp(114) <= M1(4) and M2(18);
	pp(115) <= M1(4) and M2(19);
	pp(116) <= M1(4) and M2(20);
	pp(117) <= M1(4) and M2(21);
	pp(118) <= M1(4) and M2(22);
	pp(119) <= M1(4) and M2(23);
	pp(120) <= M1(5) and M2(0);
	pp(121) <= M1(5) and M2(1);
	pp(122) <= M1(5) and M2(2);
	pp(123) <= M1(5) and M2(3);
	pp(124) <= M1(5) and M2(4);
	pp(125) <= M1(5) and M2(5);
	pp(126) <= M1(5) and M2(6);
	pp(127) <= M1(5) and M2(7);
	pp(128) <= M1(5) and M2(8);
	pp(129) <= M1(5) and M2(9);
	pp(130) <= M1(5) and M2(10);
	pp(131) <= M1(5) and M2(11);
	pp(132) <= M1(5) and M2(12);
	pp(133) <= M1(5) and M2(13);
	pp(134) <= M1(5) and M2(14);
	pp(135) <= M1(5) and M2(15);
	pp(136) <= M1(5) and M2(16);
	pp(137) <= M1(5) and M2(17);
	pp(138) <= M1(5) and M2(18);
	pp(139) <= M1(5) and M2(19);
	pp(140) <= M1(5) and M2(20);
	pp(141) <= M1(5) and M2(21);
	pp(142) <= M1(5) and M2(22);
	pp(143) <= M1(5) and M2(23);
	pp(144) <= M1(6) and M2(0);
	pp(145) <= M1(6) and M2(1);
	pp(146) <= M1(6) and M2(2);
	pp(147) <= M1(6) and M2(3);
	pp(148) <= M1(6) and M2(4);
	pp(149) <= M1(6) and M2(5);
	pp(150) <= M1(6) and M2(6);
	pp(151) <= M1(6) and M2(7);
	pp(152) <= M1(6) and M2(8);
	pp(153) <= M1(6) and M2(9);
	pp(154) <= M1(6) and M2(10);
	pp(155) <= M1(6) and M2(11);
	pp(156) <= M1(6) and M2(12);
	pp(157) <= M1(6) and M2(13);
	pp(158) <= M1(6) and M2(14);
	pp(159) <= M1(6) and M2(15);
	pp(160) <= M1(6) and M2(16);
	pp(161) <= M1(6) and M2(17);
	pp(162) <= M1(6) and M2(18);
	pp(163) <= M1(6) and M2(19);
	pp(164) <= M1(6) and M2(20);
	pp(165) <= M1(6) and M2(21);
	pp(166) <= M1(6) and M2(22);
	pp(167) <= M1(6) and M2(23);
	pp(168) <= M1(7) and M2(0);
	pp(169) <= M1(7) and M2(1);
	pp(170) <= M1(7) and M2(2);
	pp(171) <= M1(7) and M2(3);
	pp(172) <= M1(7) and M2(4);
	pp(173) <= M1(7) and M2(5);
	pp(174) <= M1(7) and M2(6);
	pp(175) <= M1(7) and M2(7);
	pp(176) <= M1(7) and M2(8);
	pp(177) <= M1(7) and M2(9);
	pp(178) <= M1(7) and M2(10);
	pp(179) <= M1(7) and M2(11);
	pp(180) <= M1(7) and M2(12);
	pp(181) <= M1(7) and M2(13);
	pp(182) <= M1(7) and M2(14);
	pp(183) <= M1(7) and M2(15);
	pp(184) <= M1(7) and M2(16);
	pp(185) <= M1(7) and M2(17);
	pp(186) <= M1(7) and M2(18);
	pp(187) <= M1(7) and M2(19);
	pp(188) <= M1(7) and M2(20);
	pp(189) <= M1(7) and M2(21);
	pp(190) <= M1(7) and M2(22);
	pp(191) <= M1(7) and M2(23);
	pp(192) <= M1(8) and M2(0);
	pp(193) <= M1(8) and M2(1);
	pp(194) <= M1(8) and M2(2);
	pp(195) <= M1(8) and M2(3);
	pp(196) <= M1(8) and M2(4);
	pp(197) <= M1(8) and M2(5);
	pp(198) <= M1(8) and M2(6);
	pp(199) <= M1(8) and M2(7);
	pp(200) <= M1(8) and M2(8);
	pp(201) <= M1(8) and M2(9);
	pp(202) <= M1(8) and M2(10);
	pp(203) <= M1(8) and M2(11);
	pp(204) <= M1(8) and M2(12);
	pp(205) <= M1(8) and M2(13);
	pp(206) <= M1(8) and M2(14);
	pp(207) <= M1(8) and M2(15);
	pp(208) <= M1(8) and M2(16);
	pp(209) <= M1(8) and M2(17);
	pp(210) <= M1(8) and M2(18);
	pp(211) <= M1(8) and M2(19);
	pp(212) <= M1(8) and M2(20);
	pp(213) <= M1(8) and M2(21);
	pp(214) <= M1(8) and M2(22);
	pp(215) <= M1(8) and M2(23);
	pp(216) <= M1(9) and M2(0);
	pp(217) <= M1(9) and M2(1);
	pp(218) <= M1(9) and M2(2);
	pp(219) <= M1(9) and M2(3);
	pp(220) <= M1(9) and M2(4);
	pp(221) <= M1(9) and M2(5);
	pp(222) <= M1(9) and M2(6);
	pp(223) <= M1(9) and M2(7);
	pp(224) <= M1(9) and M2(8);
	pp(225) <= M1(9) and M2(9);
	pp(226) <= M1(9) and M2(10);
	pp(227) <= M1(9) and M2(11);
	pp(228) <= M1(9) and M2(12);
	pp(229) <= M1(9) and M2(13);
	pp(230) <= M1(9) and M2(14);
	pp(231) <= M1(9) and M2(15);
	pp(232) <= M1(9) and M2(16);
	pp(233) <= M1(9) and M2(17);
	pp(234) <= M1(9) and M2(18);
	pp(235) <= M1(9) and M2(19);
	pp(236) <= M1(9) and M2(20);
	pp(237) <= M1(9) and M2(21);
	pp(238) <= M1(9) and M2(22);
	pp(239) <= M1(9) and M2(23);
	pp(240) <= M1(10) and M2(0);
	pp(241) <= M1(10) and M2(1);
	pp(242) <= M1(10) and M2(2);
	pp(243) <= M1(10) and M2(3);
	pp(244) <= M1(10) and M2(4);
	pp(245) <= M1(10) and M2(5);
	pp(246) <= M1(10) and M2(6);
	pp(247) <= M1(10) and M2(7);
	pp(248) <= M1(10) and M2(8);
	pp(249) <= M1(10) and M2(9);
	pp(250) <= M1(10) and M2(10);
	pp(251) <= M1(10) and M2(11);
	pp(252) <= M1(10) and M2(12);
	pp(253) <= M1(10) and M2(13);
	pp(254) <= M1(10) and M2(14);
	pp(255) <= M1(10) and M2(15);
	pp(256) <= M1(10) and M2(16);
	pp(257) <= M1(10) and M2(17);
	pp(258) <= M1(10) and M2(18);
	pp(259) <= M1(10) and M2(19);
	pp(260) <= M1(10) and M2(20);
	pp(261) <= M1(10) and M2(21);
	pp(262) <= M1(10) and M2(22);
	pp(263) <= M1(10) and M2(23);
	pp(264) <= M1(11) and M2(0);
	pp(265) <= M1(11) and M2(1);
	pp(266) <= M1(11) and M2(2);
	pp(267) <= M1(11) and M2(3);
	pp(268) <= M1(11) and M2(4);
	pp(269) <= M1(11) and M2(5);
	pp(270) <= M1(11) and M2(6);
	pp(271) <= M1(11) and M2(7);
	pp(272) <= M1(11) and M2(8);
	pp(273) <= M1(11) and M2(9);
	pp(274) <= M1(11) and M2(10);
	pp(275) <= M1(11) and M2(11);
	pp(276) <= M1(11) and M2(12);
	pp(277) <= M1(11) and M2(13);
	pp(278) <= M1(11) and M2(14);
	pp(279) <= M1(11) and M2(15);
	pp(280) <= M1(11) and M2(16);
	pp(281) <= M1(11) and M2(17);
	pp(282) <= M1(11) and M2(18);
	pp(283) <= M1(11) and M2(19);
	pp(284) <= M1(11) and M2(20);
	pp(285) <= M1(11) and M2(21);
	pp(286) <= M1(11) and M2(22);
	pp(287) <= M1(11) and M2(23);
	pp(288) <= M1(12) and M2(0);
	pp(289) <= M1(12) and M2(1);
	pp(290) <= M1(12) and M2(2);
	pp(291) <= M1(12) and M2(3);
	pp(292) <= M1(12) and M2(4);
	pp(293) <= M1(12) and M2(5);
	pp(294) <= M1(12) and M2(6);
	pp(295) <= M1(12) and M2(7);
	pp(296) <= M1(12) and M2(8);
	pp(297) <= M1(12) and M2(9);
	pp(298) <= M1(12) and M2(10);
	pp(299) <= M1(12) and M2(11);
	pp(300) <= M1(12) and M2(12);
	pp(301) <= M1(12) and M2(13);
	pp(302) <= M1(12) and M2(14);
	pp(303) <= M1(12) and M2(15);
	pp(304) <= M1(12) and M2(16);
	pp(305) <= M1(12) and M2(17);
	pp(306) <= M1(12) and M2(18);
	pp(307) <= M1(12) and M2(19);
	pp(308) <= M1(12) and M2(20);
	pp(309) <= M1(12) and M2(21);
	pp(310) <= M1(12) and M2(22);
	pp(311) <= M1(12) and M2(23);
	pp(312) <= M1(13) and M2(0);
	pp(313) <= M1(13) and M2(1);
	pp(314) <= M1(13) and M2(2);
	pp(315) <= M1(13) and M2(3);
	pp(316) <= M1(13) and M2(4);
	pp(317) <= M1(13) and M2(5);
	pp(318) <= M1(13) and M2(6);
	pp(319) <= M1(13) and M2(7);
	pp(320) <= M1(13) and M2(8);
	pp(321) <= M1(13) and M2(9);
	pp(322) <= M1(13) and M2(10);
	pp(323) <= M1(13) and M2(11);
	pp(324) <= M1(13) and M2(12);
	pp(325) <= M1(13) and M2(13);
	pp(326) <= M1(13) and M2(14);
	pp(327) <= M1(13) and M2(15);
	pp(328) <= M1(13) and M2(16);
	pp(329) <= M1(13) and M2(17);
	pp(330) <= M1(13) and M2(18);
	pp(331) <= M1(13) and M2(19);
	pp(332) <= M1(13) and M2(20);
	pp(333) <= M1(13) and M2(21);
	pp(334) <= M1(13) and M2(22);
	pp(335) <= M1(13) and M2(23);
	pp(336) <= M1(14) and M2(0);
	pp(337) <= M1(14) and M2(1);
	pp(338) <= M1(14) and M2(2);
	pp(339) <= M1(14) and M2(3);
	pp(340) <= M1(14) and M2(4);
	pp(341) <= M1(14) and M2(5);
	pp(342) <= M1(14) and M2(6);
	pp(343) <= M1(14) and M2(7);
	pp(344) <= M1(14) and M2(8);
	pp(345) <= M1(14) and M2(9);
	pp(346) <= M1(14) and M2(10);
	pp(347) <= M1(14) and M2(11);
	pp(348) <= M1(14) and M2(12);
	pp(349) <= M1(14) and M2(13);
	pp(350) <= M1(14) and M2(14);
	pp(351) <= M1(14) and M2(15);
	pp(352) <= M1(14) and M2(16);
	pp(353) <= M1(14) and M2(17);
	pp(354) <= M1(14) and M2(18);
	pp(355) <= M1(14) and M2(19);
	pp(356) <= M1(14) and M2(20);
	pp(357) <= M1(14) and M2(21);
	pp(358) <= M1(14) and M2(22);
	pp(359) <= M1(14) and M2(23);
	pp(360) <= M1(15) and M2(0);
	pp(361) <= M1(15) and M2(1);
	pp(362) <= M1(15) and M2(2);
	pp(363) <= M1(15) and M2(3);
	pp(364) <= M1(15) and M2(4);
	pp(365) <= M1(15) and M2(5);
	pp(366) <= M1(15) and M2(6);
	pp(367) <= M1(15) and M2(7);
	pp(368) <= M1(15) and M2(8);
	pp(369) <= M1(15) and M2(9);
	pp(370) <= M1(15) and M2(10);
	pp(371) <= M1(15) and M2(11);
	pp(372) <= M1(15) and M2(12);
	pp(373) <= M1(15) and M2(13);
	pp(374) <= M1(15) and M2(14);
	pp(375) <= M1(15) and M2(15);
	pp(376) <= M1(15) and M2(16);
	pp(377) <= M1(15) and M2(17);
	pp(378) <= M1(15) and M2(18);
	pp(379) <= M1(15) and M2(19);
	pp(380) <= M1(15) and M2(20);
	pp(381) <= M1(15) and M2(21);
	pp(382) <= M1(15) and M2(22);
	pp(383) <= M1(15) and M2(23);
	pp(384) <= M1(16) and M2(0);
	pp(385) <= M1(16) and M2(1);
	pp(386) <= M1(16) and M2(2);
	pp(387) <= M1(16) and M2(3);
	pp(388) <= M1(16) and M2(4);
	pp(389) <= M1(16) and M2(5);
	pp(390) <= M1(16) and M2(6);
	pp(391) <= M1(16) and M2(7);
	pp(392) <= M1(16) and M2(8);
	pp(393) <= M1(16) and M2(9);
	pp(394) <= M1(16) and M2(10);
	pp(395) <= M1(16) and M2(11);
	pp(396) <= M1(16) and M2(12);
	pp(397) <= M1(16) and M2(13);
	pp(398) <= M1(16) and M2(14);
	pp(399) <= M1(16) and M2(15);
	pp(400) <= M1(16) and M2(16);
	pp(401) <= M1(16) and M2(17);
	pp(402) <= M1(16) and M2(18);
	pp(403) <= M1(16) and M2(19);
	pp(404) <= M1(16) and M2(20);
	pp(405) <= M1(16) and M2(21);
	pp(406) <= M1(16) and M2(22);
	pp(407) <= M1(16) and M2(23);
	pp(408) <= M1(17) and M2(0);
	pp(409) <= M1(17) and M2(1);
	pp(410) <= M1(17) and M2(2);
	pp(411) <= M1(17) and M2(3);
	pp(412) <= M1(17) and M2(4);
	pp(413) <= M1(17) and M2(5);
	pp(414) <= M1(17) and M2(6);
	pp(415) <= M1(17) and M2(7);
	pp(416) <= M1(17) and M2(8);
	pp(417) <= M1(17) and M2(9);
	pp(418) <= M1(17) and M2(10);
	pp(419) <= M1(17) and M2(11);
	pp(420) <= M1(17) and M2(12);
	pp(421) <= M1(17) and M2(13);
	pp(422) <= M1(17) and M2(14);
	pp(423) <= M1(17) and M2(15);
	pp(424) <= M1(17) and M2(16);
	pp(425) <= M1(17) and M2(17);
	pp(426) <= M1(17) and M2(18);
	pp(427) <= M1(17) and M2(19);
	pp(428) <= M1(17) and M2(20);
	pp(429) <= M1(17) and M2(21);
	pp(430) <= M1(17) and M2(22);
	pp(431) <= M1(17) and M2(23);
	pp(432) <= M1(18) and M2(0);
	pp(433) <= M1(18) and M2(1);
	pp(434) <= M1(18) and M2(2);
	pp(435) <= M1(18) and M2(3);
	pp(436) <= M1(18) and M2(4);
	pp(437) <= M1(18) and M2(5);
	pp(438) <= M1(18) and M2(6);
	pp(439) <= M1(18) and M2(7);
	pp(440) <= M1(18) and M2(8);
	pp(441) <= M1(18) and M2(9);
	pp(442) <= M1(18) and M2(10);
	pp(443) <= M1(18) and M2(11);
	pp(444) <= M1(18) and M2(12);
	pp(445) <= M1(18) and M2(13);
	pp(446) <= M1(18) and M2(14);
	pp(447) <= M1(18) and M2(15);
	pp(448) <= M1(18) and M2(16);
	pp(449) <= M1(18) and M2(17);
	pp(450) <= M1(18) and M2(18);
	pp(451) <= M1(18) and M2(19);
	pp(452) <= M1(18) and M2(20);
	pp(453) <= M1(18) and M2(21);
	pp(454) <= M1(18) and M2(22);
	pp(455) <= M1(18) and M2(23);
	pp(456) <= M1(19) and M2(0);
	pp(457) <= M1(19) and M2(1);
	pp(458) <= M1(19) and M2(2);
	pp(459) <= M1(19) and M2(3);
	pp(460) <= M1(19) and M2(4);
	pp(461) <= M1(19) and M2(5);
	pp(462) <= M1(19) and M2(6);
	pp(463) <= M1(19) and M2(7);
	pp(464) <= M1(19) and M2(8);
	pp(465) <= M1(19) and M2(9);
	pp(466) <= M1(19) and M2(10);
	pp(467) <= M1(19) and M2(11);
	pp(468) <= M1(19) and M2(12);
	pp(469) <= M1(19) and M2(13);
	pp(470) <= M1(19) and M2(14);
	pp(471) <= M1(19) and M2(15);
	pp(472) <= M1(19) and M2(16);
	pp(473) <= M1(19) and M2(17);
	pp(474) <= M1(19) and M2(18);
	pp(475) <= M1(19) and M2(19);
	pp(476) <= M1(19) and M2(20);
	pp(477) <= M1(19) and M2(21);
	pp(478) <= M1(19) and M2(22);
	pp(479) <= M1(19) and M2(23);
	pp(480) <= M1(20) and M2(0);
	pp(481) <= M1(20) and M2(1);
	pp(482) <= M1(20) and M2(2);
	pp(483) <= M1(20) and M2(3);
	pp(484) <= M1(20) and M2(4);
	pp(485) <= M1(20) and M2(5);
	pp(486) <= M1(20) and M2(6);
	pp(487) <= M1(20) and M2(7);
	pp(488) <= M1(20) and M2(8);
	pp(489) <= M1(20) and M2(9);
	pp(490) <= M1(20) and M2(10);
	pp(491) <= M1(20) and M2(11);
	pp(492) <= M1(20) and M2(12);
	pp(493) <= M1(20) and M2(13);
	pp(494) <= M1(20) and M2(14);
	pp(495) <= M1(20) and M2(15);
	pp(496) <= M1(20) and M2(16);
	pp(497) <= M1(20) and M2(17);
	pp(498) <= M1(20) and M2(18);
	pp(499) <= M1(20) and M2(19);
	pp(500) <= M1(20) and M2(20);
	pp(501) <= M1(20) and M2(21);
	pp(502) <= M1(20) and M2(22);
	pp(503) <= M1(20) and M2(23);
	pp(504) <= M1(21) and M2(0);
	pp(505) <= M1(21) and M2(1);
	pp(506) <= M1(21) and M2(2);
	pp(507) <= M1(21) and M2(3);
	pp(508) <= M1(21) and M2(4);
	pp(509) <= M1(21) and M2(5);
	pp(510) <= M1(21) and M2(6);
	pp(511) <= M1(21) and M2(7);
	pp(512) <= M1(21) and M2(8);
	pp(513) <= M1(21) and M2(9);
	pp(514) <= M1(21) and M2(10);
	pp(515) <= M1(21) and M2(11);
	pp(516) <= M1(21) and M2(12);
	pp(517) <= M1(21) and M2(13);
	pp(518) <= M1(21) and M2(14);
	pp(519) <= M1(21) and M2(15);
	pp(520) <= M1(21) and M2(16);
	pp(521) <= M1(21) and M2(17);
	pp(522) <= M1(21) and M2(18);
	pp(523) <= M1(21) and M2(19);
	pp(524) <= M1(21) and M2(20);
	pp(525) <= M1(21) and M2(21);
	pp(526) <= M1(21) and M2(22);
	pp(527) <= M1(21) and M2(23);
	pp(528) <= M1(22) and M2(0);
	pp(529) <= M1(22) and M2(1);
	pp(530) <= M1(22) and M2(2);
	pp(531) <= M1(22) and M2(3);
	pp(532) <= M1(22) and M2(4);
	pp(533) <= M1(22) and M2(5);
	pp(534) <= M1(22) and M2(6);
	pp(535) <= M1(22) and M2(7);
	pp(536) <= M1(22) and M2(8);
	pp(537) <= M1(22) and M2(9);
	pp(538) <= M1(22) and M2(10);
	pp(539) <= M1(22) and M2(11);
	pp(540) <= M1(22) and M2(12);
	pp(541) <= M1(22) and M2(13);
	pp(542) <= M1(22) and M2(14);
	pp(543) <= M1(22) and M2(15);
	pp(544) <= M1(22) and M2(16);
	pp(545) <= M1(22) and M2(17);
	pp(546) <= M1(22) and M2(18);
	pp(547) <= M1(22) and M2(19);
	pp(548) <= M1(22) and M2(20);
	pp(549) <= M1(22) and M2(21);
	pp(550) <= M1(22) and M2(22);
	pp(551) <= M1(22) and M2(23);
	pp(552) <= M1(23) and M2(0);
	pp(553) <= M1(23) and M2(1);
	pp(554) <= M1(23) and M2(2);
	pp(555) <= M1(23) and M2(3);
	pp(556) <= M1(23) and M2(4);
	pp(557) <= M1(23) and M2(5);
	pp(558) <= M1(23) and M2(6);
	pp(559) <= M1(23) and M2(7);
	pp(560) <= M1(23) and M2(8);
	pp(561) <= M1(23) and M2(9);
	pp(562) <= M1(23) and M2(10);
	pp(563) <= M1(23) and M2(11);
	pp(564) <= M1(23) and M2(12);
	pp(565) <= M1(23) and M2(13);
	pp(566) <= M1(23) and M2(14);
	pp(567) <= M1(23) and M2(15);
	pp(568) <= M1(23) and M2(16);
	pp(569) <= M1(23) and M2(17);
	pp(570) <= M1(23) and M2(18);
	pp(571) <= M1(23) and M2(19);
	pp(572) <= M1(23) and M2(20);
	pp(573) <= M1(23) and M2(21);
	pp(574) <= M1(23) and M2(22);
	pp(575) <= M1(23) and M2(23);
	

	-- ALLOCATE ADDERS
	-- Stage J = 7; d_7 = 19
	-- HAs ALLOCATED: 6 (6 TOTAL)
	-- FAs ALLOCATED: 24 (24 TOTAL)
	HA_1: HA port map(pp(456), pp(433), sum(0), carry(0));
	FA_2: FA port map(pp(480), pp(457), pp(434), sum(1), carry(1));
	HA_3: HA port map(pp(411), pp(388), sum(2), carry(2));
	FA_4: FA port map(pp(504), pp(481), pp(458), sum(3), carry(3));
	FA_5: FA port map(pp(435), pp(412), pp(389), sum(4), carry(4));
	HA_6: HA port map(pp(366), pp(343), sum(5), carry(5));
	FA_7: FA port map(pp(528), pp(505), pp(482), sum(6), carry(6));
	FA_8: FA port map(pp(459), pp(436), pp(413), sum(7), carry(7));
	FA_9: FA port map(pp(390), pp(367), pp(344), sum(8), carry(8));
	HA_10: HA port map(pp(321), pp(298), sum(9), carry(9));
	FA_11: FA port map(pp(552), pp(529), pp(506), sum(10), carry(10));
	FA_12: FA port map(pp(483), pp(460), pp(437), sum(11), carry(11));
	FA_13: FA port map(pp(414), pp(391), pp(368), sum(12), carry(12));
	FA_14: FA port map(pp(345), pp(322), pp(299), sum(13), carry(13));
	HA_15: HA port map(pp(276), pp(253), sum(14), carry(14));
	FA_16: FA port map(pp(553), pp(530), pp(507), sum(15), carry(15));
	FA_17: FA port map(pp(484), pp(461), pp(438), sum(16), carry(16));
	FA_18: FA port map(pp(415), pp(392), pp(369), sum(17), carry(17));
	FA_19: FA port map(pp(346), pp(323), pp(300), sum(18), carry(18));
	HA_20: HA port map(pp(277), pp(254), sum(19), carry(19));
	FA_21: FA port map(pp(554), pp(531), pp(508), sum(20), carry(20));
	FA_22: FA port map(pp(485), pp(462), pp(439), sum(21), carry(21));
	FA_23: FA port map(pp(416), pp(393), pp(370), sum(22), carry(22));
	FA_24: FA port map(pp(347), pp(324), pp(301), sum(23), carry(23));
	FA_25: FA port map(pp(555), pp(532), pp(509), sum(24), carry(24));
	FA_26: FA port map(pp(486), pp(463), pp(440), sum(25), carry(25));
	FA_27: FA port map(pp(417), pp(394), pp(371), sum(26), carry(26));
	FA_28: FA port map(pp(556), pp(533), pp(510), sum(27), carry(27));
	FA_29: FA port map(pp(487), pp(464), pp(441), sum(28), carry(28));
	FA_30: FA port map(pp(557), pp(534), pp(511), sum(29), carry(29));
	
	-- Stage J = 6; d_6 = 13
	-- HAs ALLOCATED: 6 (12 TOTAL)
	-- FAs ALLOCATED: 96 (120 TOTAL)
	HA_31: HA port map(pp(312), pp(289), sum(30), carry(30));
	FA_32: FA port map(pp(336), pp(313), pp(290), sum(31), carry(31));
	HA_33: HA port map(pp(267), pp(244), sum(32), carry(32));
	FA_34: FA port map(pp(360), pp(337), pp(314), sum(33), carry(33));
	FA_35: FA port map(pp(291), pp(268), pp(245), sum(34), carry(34));
	HA_36: HA port map(pp(222), pp(199), sum(35), carry(35));
	FA_37: FA port map(pp(384), pp(361), pp(338), sum(36), carry(36));
	FA_38: FA port map(pp(315), pp(292), pp(269), sum(37), carry(37));
	FA_39: FA port map(pp(246), pp(223), pp(200), sum(38), carry(38));
	HA_40: HA port map(pp(177), pp(154), sum(39), carry(39));
	FA_41: FA port map(pp(408), pp(385), pp(362), sum(40), carry(40));
	FA_42: FA port map(pp(339), pp(316), pp(293), sum(41), carry(41));
	FA_43: FA port map(pp(270), pp(247), pp(224), sum(42), carry(42));
	FA_44: FA port map(pp(201), pp(178), pp(155), sum(43), carry(43));
	HA_45: HA port map(pp(132), pp(109), sum(44), carry(44));
	FA_46: FA port map(pp(432), pp(409), pp(386), sum(45), carry(45));
	FA_47: FA port map(pp(363), pp(340), pp(317), sum(46), carry(46));
	FA_48: FA port map(pp(294), pp(271), pp(248), sum(47), carry(47));
	FA_49: FA port map(pp(225), pp(202), pp(179), sum(48), carry(48));
	FA_50: FA port map(pp(156), pp(133), pp(110), sum(49), carry(49));
	HA_51: HA port map(pp(87), pp(64), sum(50), carry(50));
	FA_52: FA port map(pp(410), pp(387), pp(364), sum(51), carry(51));
	FA_53: FA port map(pp(341), pp(318), pp(295), sum(52), carry(52));
	FA_54: FA port map(pp(272), pp(249), pp(226), sum(53), carry(53));
	FA_55: FA port map(pp(203), pp(180), pp(157), sum(54), carry(54));
	FA_56: FA port map(pp(134), pp(111), pp(88), sum(55), carry(55));
	FA_57: FA port map(pp(65), pp(42), pp(19), sum(56), carry(56));
	FA_58: FA port map(pp(365), pp(342), pp(319), sum(57), carry(57));
	FA_59: FA port map(pp(296), pp(273), pp(250), sum(58), carry(58));
	FA_60: FA port map(pp(227), pp(204), pp(181), sum(59), carry(59));
	FA_61: FA port map(pp(158), pp(135), pp(112), sum(60), carry(60));
	FA_62: FA port map(pp(89), pp(66), pp(43), sum(61), carry(61));
	FA_63: FA port map(pp(20), carry(0), sum(1), sum(62), carry(62));
	FA_64: FA port map(pp(320), pp(297), pp(274), sum(63), carry(63));
	FA_65: FA port map(pp(251), pp(228), pp(205), sum(64), carry(64));
	FA_66: FA port map(pp(182), pp(159), pp(136), sum(65), carry(65));
	FA_67: FA port map(pp(113), pp(90), pp(67), sum(66), carry(66));
	FA_68: FA port map(pp(44), pp(21), carry(2), sum(67), carry(67));
	FA_69: FA port map(carry(1), sum(3), sum(4), sum(68), carry(68));
	FA_70: FA port map(pp(275), pp(252), pp(229), sum(69), carry(69));
	FA_71: FA port map(pp(206), pp(183), pp(160), sum(70), carry(70));
	FA_72: FA port map(pp(137), pp(114), pp(91), sum(71), carry(71));
	FA_73: FA port map(pp(68), pp(45), pp(22), sum(72), carry(72));
	FA_74: FA port map(carry(5), carry(4), carry(3), sum(73), carry(73));
	FA_75: FA port map(sum(6), sum(7), sum(8), sum(74), carry(74));
	FA_76: FA port map(pp(230), pp(207), pp(184), sum(75), carry(75));
	FA_77: FA port map(pp(161), pp(138), pp(115), sum(76), carry(76));
	FA_78: FA port map(pp(92), pp(69), pp(46), sum(77), carry(77));
	FA_79: FA port map(pp(23), carry(9), carry(8), sum(78), carry(78));
	FA_80: FA port map(carry(7), carry(6), sum(10), sum(79), carry(79));
	FA_81: FA port map(sum(11), sum(12), sum(13), sum(80), carry(80));
	FA_82: FA port map(pp(231), pp(208), pp(185), sum(81), carry(81));
	FA_83: FA port map(pp(162), pp(139), pp(116), sum(82), carry(82));
	FA_84: FA port map(pp(93), pp(70), pp(47), sum(83), carry(83));
	FA_85: FA port map(carry(14), carry(13), carry(12), sum(84), carry(84));
	FA_86: FA port map(carry(11), carry(10), sum(15), sum(85), carry(85));
	FA_87: FA port map(sum(16), sum(17), sum(18), sum(86), carry(86));
	FA_88: FA port map(pp(278), pp(255), pp(232), sum(87), carry(87));
	FA_89: FA port map(pp(209), pp(186), pp(163), sum(88), carry(88));
	FA_90: FA port map(pp(140), pp(117), pp(94), sum(89), carry(89));
	FA_91: FA port map(pp(71), carry(19), carry(18), sum(90), carry(90));
	FA_92: FA port map(carry(17), carry(16), carry(15), sum(91), carry(91));
	FA_93: FA port map(sum(20), sum(21), sum(22), sum(92), carry(92));
	FA_94: FA port map(pp(348), pp(325), pp(302), sum(93), carry(93));
	FA_95: FA port map(pp(279), pp(256), pp(233), sum(94), carry(94));
	FA_96: FA port map(pp(210), pp(187), pp(164), sum(95), carry(95));
	FA_97: FA port map(pp(141), pp(118), pp(95), sum(96), carry(96));
	FA_98: FA port map(carry(23), carry(22), carry(21), sum(97), carry(97));
	FA_99: FA port map(carry(20), sum(24), sum(25), sum(98), carry(98));
	FA_100: FA port map(pp(418), pp(395), pp(372), sum(99), carry(99));
	FA_101: FA port map(pp(349), pp(326), pp(303), sum(100), carry(100));
	FA_102: FA port map(pp(280), pp(257), pp(234), sum(101), carry(101));
	FA_103: FA port map(pp(211), pp(188), pp(165), sum(102), carry(102));
	FA_104: FA port map(pp(142), pp(119), carry(26), sum(103), carry(103));
	FA_105: FA port map(carry(25), carry(24), sum(27), sum(104), carry(104));
	FA_106: FA port map(pp(488), pp(465), pp(442), sum(105), carry(105));
	FA_107: FA port map(pp(419), pp(396), pp(373), sum(106), carry(106));
	FA_108: FA port map(pp(350), pp(327), pp(304), sum(107), carry(107));
	FA_109: FA port map(pp(281), pp(258), pp(235), sum(108), carry(108));
	FA_110: FA port map(pp(212), pp(189), pp(166), sum(109), carry(109));
	FA_111: FA port map(pp(143), carry(28), carry(27), sum(110), carry(110));
	FA_112: FA port map(pp(558), pp(535), pp(512), sum(111), carry(111));
	FA_113: FA port map(pp(489), pp(466), pp(443), sum(112), carry(112));
	FA_114: FA port map(pp(420), pp(397), pp(374), sum(113), carry(113));
	FA_115: FA port map(pp(351), pp(328), pp(305), sum(114), carry(114));
	FA_116: FA port map(pp(282), pp(259), pp(236), sum(115), carry(115));
	FA_117: FA port map(pp(213), pp(190), pp(167), sum(116), carry(116));
	FA_118: FA port map(pp(559), pp(536), pp(513), sum(117), carry(117));
	FA_119: FA port map(pp(490), pp(467), pp(444), sum(118), carry(118));
	FA_120: FA port map(pp(421), pp(398), pp(375), sum(119), carry(119));
	FA_121: FA port map(pp(352), pp(329), pp(306), sum(120), carry(120));
	FA_122: FA port map(pp(283), pp(260), pp(237), sum(121), carry(121));
	FA_123: FA port map(pp(560), pp(537), pp(514), sum(122), carry(122));
	FA_124: FA port map(pp(491), pp(468), pp(445), sum(123), carry(123));
	FA_125: FA port map(pp(422), pp(399), pp(376), sum(124), carry(124));
	FA_126: FA port map(pp(353), pp(330), pp(307), sum(125), carry(125));
	FA_127: FA port map(pp(561), pp(538), pp(515), sum(126), carry(126));
	FA_128: FA port map(pp(492), pp(469), pp(446), sum(127), carry(127));
	FA_129: FA port map(pp(423), pp(400), pp(377), sum(128), carry(128));
	FA_130: FA port map(pp(562), pp(539), pp(516), sum(129), carry(129));
	FA_131: FA port map(pp(493), pp(470), pp(447), sum(130), carry(130));
	FA_132: FA port map(pp(563), pp(540), pp(517), sum(131), carry(131));
	
	-- Stage J = 5; d_5 = 9
	-- HAs ALLOCATED: 4 (16 TOTAL)
	-- FAs ALLOCATED: 104 (224 TOTAL)
	HA_133: HA port map(pp(216), pp(193), sum(132), carry(132));
	FA_134: FA port map(pp(240), pp(217), pp(194), sum(133), carry(133));
	HA_135: HA port map(pp(171), pp(148), sum(134), carry(134));
	FA_136: FA port map(pp(264), pp(241), pp(218), sum(135), carry(135));
	FA_137: FA port map(pp(195), pp(172), pp(149), sum(136), carry(136));
	HA_138: HA port map(pp(126), pp(103), sum(137), carry(137));
	FA_139: FA port map(pp(288), pp(265), pp(242), sum(138), carry(138));
	FA_140: FA port map(pp(219), pp(196), pp(173), sum(139), carry(139));
	FA_141: FA port map(pp(150), pp(127), pp(104), sum(140), carry(140));
	HA_142: HA port map(pp(81), pp(58), sum(141), carry(141));
	FA_143: FA port map(pp(266), pp(243), pp(220), sum(142), carry(142));
	FA_144: FA port map(pp(197), pp(174), pp(151), sum(143), carry(143));
	FA_145: FA port map(pp(128), pp(105), pp(82), sum(144), carry(144));
	FA_146: FA port map(pp(59), pp(36), pp(13), sum(145), carry(145));
	FA_147: FA port map(pp(221), pp(198), pp(175), sum(146), carry(146));
	FA_148: FA port map(pp(152), pp(129), pp(106), sum(147), carry(147));
	FA_149: FA port map(pp(83), pp(60), pp(37), sum(148), carry(148));
	FA_150: FA port map(pp(14), carry(30), sum(31), sum(149), carry(149));
	FA_151: FA port map(pp(176), pp(153), pp(130), sum(150), carry(150));
	FA_152: FA port map(pp(107), pp(84), pp(61), sum(151), carry(151));
	FA_153: FA port map(pp(38), pp(15), carry(32), sum(152), carry(152));
	FA_154: FA port map(carry(31), sum(33), sum(34), sum(153), carry(153));
	FA_155: FA port map(pp(131), pp(108), pp(85), sum(154), carry(154));
	FA_156: FA port map(pp(62), pp(39), pp(16), sum(155), carry(155));
	FA_157: FA port map(carry(35), carry(34), carry(33), sum(156), carry(156));
	FA_158: FA port map(sum(36), sum(37), sum(38), sum(157), carry(157));
	FA_159: FA port map(pp(86), pp(63), pp(40), sum(158), carry(158));
	FA_160: FA port map(pp(17), carry(39), carry(38), sum(159), carry(159));
	FA_161: FA port map(carry(37), carry(36), sum(40), sum(160), carry(160));
	FA_162: FA port map(sum(41), sum(42), sum(43), sum(161), carry(161));
	FA_163: FA port map(pp(41), pp(18), carry(44), sum(162), carry(162));
	FA_164: FA port map(carry(43), carry(42), carry(41), sum(163), carry(163));
	FA_165: FA port map(carry(40), sum(45), sum(46), sum(164), carry(164));
	FA_166: FA port map(sum(47), sum(48), sum(49), sum(165), carry(165));
	FA_167: FA port map(sum(0), carry(50), carry(49), sum(166), carry(166));
	FA_168: FA port map(carry(48), carry(47), carry(46), sum(167), carry(167));
	FA_169: FA port map(carry(45), sum(51), sum(52), sum(168), carry(168));
	FA_170: FA port map(sum(53), sum(54), sum(55), sum(169), carry(169));
	FA_171: FA port map(sum(2), carry(56), carry(55), sum(170), carry(170));
	FA_172: FA port map(carry(54), carry(53), carry(52), sum(171), carry(171));
	FA_173: FA port map(carry(51), sum(57), sum(58), sum(172), carry(172));
	FA_174: FA port map(sum(59), sum(60), sum(61), sum(173), carry(173));
	FA_175: FA port map(sum(5), carry(62), carry(61), sum(174), carry(174));
	FA_176: FA port map(carry(60), carry(59), carry(58), sum(175), carry(175));
	FA_177: FA port map(carry(57), sum(63), sum(64), sum(176), carry(176));
	FA_178: FA port map(sum(65), sum(66), sum(67), sum(177), carry(177));
	FA_179: FA port map(sum(9), carry(68), carry(67), sum(178), carry(178));
	FA_180: FA port map(carry(66), carry(65), carry(64), sum(179), carry(179));
	FA_181: FA port map(carry(63), sum(69), sum(70), sum(180), carry(180));
	FA_182: FA port map(sum(71), sum(72), sum(73), sum(181), carry(181));
	FA_183: FA port map(sum(14), carry(74), carry(73), sum(182), carry(182));
	FA_184: FA port map(carry(72), carry(71), carry(70), sum(183), carry(183));
	FA_185: FA port map(carry(69), sum(75), sum(76), sum(184), carry(184));
	FA_186: FA port map(sum(77), sum(78), sum(79), sum(185), carry(185));
	FA_187: FA port map(sum(19), carry(80), carry(79), sum(186), carry(186));
	FA_188: FA port map(carry(78), carry(77), carry(76), sum(187), carry(187));
	FA_189: FA port map(carry(75), sum(81), sum(82), sum(188), carry(188));
	FA_190: FA port map(sum(83), sum(84), sum(85), sum(189), carry(189));
	FA_191: FA port map(sum(23), carry(86), carry(85), sum(190), carry(190));
	FA_192: FA port map(carry(84), carry(83), carry(82), sum(191), carry(191));
	FA_193: FA port map(carry(81), sum(87), sum(88), sum(192), carry(192));
	FA_194: FA port map(sum(89), sum(90), sum(91), sum(193), carry(193));
	FA_195: FA port map(sum(26), carry(92), carry(91), sum(194), carry(194));
	FA_196: FA port map(carry(90), carry(89), carry(88), sum(195), carry(195));
	FA_197: FA port map(carry(87), sum(93), sum(94), sum(196), carry(196));
	FA_198: FA port map(sum(95), sum(96), sum(97), sum(197), carry(197));
	FA_199: FA port map(sum(28), carry(98), carry(97), sum(198), carry(198));
	FA_200: FA port map(carry(96), carry(95), carry(94), sum(199), carry(199));
	FA_201: FA port map(carry(93), sum(99), sum(100), sum(200), carry(200));
	FA_202: FA port map(sum(101), sum(102), sum(103), sum(201), carry(201));
	FA_203: FA port map(sum(29), carry(104), carry(103), sum(202), carry(202));
	FA_204: FA port map(carry(102), carry(101), carry(100), sum(203), carry(203));
	FA_205: FA port map(carry(99), sum(105), sum(106), sum(204), carry(204));
	FA_206: FA port map(sum(107), sum(108), sum(109), sum(205), carry(205));
	FA_207: FA port map(carry(29), carry(110), carry(109), sum(206), carry(206));
	FA_208: FA port map(carry(108), carry(107), carry(106), sum(207), carry(207));
	FA_209: FA port map(carry(105), sum(111), sum(112), sum(208), carry(208));
	FA_210: FA port map(sum(113), sum(114), sum(115), sum(209), carry(209));
	FA_211: FA port map(pp(214), pp(191), carry(116), sum(210), carry(210));
	FA_212: FA port map(carry(115), carry(114), carry(113), sum(211), carry(211));
	FA_213: FA port map(carry(112), carry(111), sum(117), sum(212), carry(212));
	FA_214: FA port map(sum(118), sum(119), sum(120), sum(213), carry(213));
	FA_215: FA port map(pp(284), pp(261), pp(238), sum(214), carry(214));
	FA_216: FA port map(pp(215), carry(121), carry(120), sum(215), carry(215));
	FA_217: FA port map(carry(119), carry(118), carry(117), sum(216), carry(216));
	FA_218: FA port map(sum(122), sum(123), sum(124), sum(217), carry(217));
	FA_219: FA port map(pp(354), pp(331), pp(308), sum(218), carry(218));
	FA_220: FA port map(pp(285), pp(262), pp(239), sum(219), carry(219));
	FA_221: FA port map(carry(125), carry(124), carry(123), sum(220), carry(220));
	FA_222: FA port map(carry(122), sum(126), sum(127), sum(221), carry(221));
	FA_223: FA port map(pp(424), pp(401), pp(378), sum(222), carry(222));
	FA_224: FA port map(pp(355), pp(332), pp(309), sum(223), carry(223));
	FA_225: FA port map(pp(286), pp(263), carry(128), sum(224), carry(224));
	FA_226: FA port map(carry(127), carry(126), sum(129), sum(225), carry(225));
	FA_227: FA port map(pp(494), pp(471), pp(448), sum(226), carry(226));
	FA_228: FA port map(pp(425), pp(402), pp(379), sum(227), carry(227));
	FA_229: FA port map(pp(356), pp(333), pp(310), sum(228), carry(228));
	FA_230: FA port map(pp(287), carry(130), carry(129), sum(229), carry(229));
	FA_231: FA port map(pp(564), pp(541), pp(518), sum(230), carry(230));
	FA_232: FA port map(pp(495), pp(472), pp(449), sum(231), carry(231));
	FA_233: FA port map(pp(426), pp(403), pp(380), sum(232), carry(232));
	FA_234: FA port map(pp(357), pp(334), pp(311), sum(233), carry(233));
	FA_235: FA port map(pp(565), pp(542), pp(519), sum(234), carry(234));
	FA_236: FA port map(pp(496), pp(473), pp(450), sum(235), carry(235));
	FA_237: FA port map(pp(427), pp(404), pp(381), sum(236), carry(236));
	FA_238: FA port map(pp(566), pp(543), pp(520), sum(237), carry(237));
	FA_239: FA port map(pp(497), pp(474), pp(451), sum(238), carry(238));
	FA_240: FA port map(pp(567), pp(544), pp(521), sum(239), carry(239));
	
	-- Stage J = 4; d_4 = 6
	-- HAs ALLOCATED: 3 (19 TOTAL)
	-- FAs ALLOCATED: 99 (323 TOTAL)
	HA_241: HA port map(pp(144), pp(121), sum(240), carry(240));
	FA_242: FA port map(pp(168), pp(145), pp(122), sum(241), carry(241));
	HA_243: HA port map(pp(99), pp(76), sum(242), carry(242));
	FA_244: FA port map(pp(192), pp(169), pp(146), sum(243), carry(243));
	FA_245: FA port map(pp(123), pp(100), pp(77), sum(244), carry(244));
	HA_246: HA port map(pp(54), pp(31), sum(245), carry(245));
	FA_247: FA port map(pp(170), pp(147), pp(124), sum(246), carry(246));
	FA_248: FA port map(pp(101), pp(78), pp(55), sum(247), carry(247));
	FA_249: FA port map(pp(32), pp(9), sum(132), sum(248), carry(248));
	FA_250: FA port map(pp(125), pp(102), pp(79), sum(249), carry(249));
	FA_251: FA port map(pp(56), pp(33), pp(10), sum(250), carry(250));
	FA_252: FA port map(carry(132), sum(133), sum(134), sum(251), carry(251));
	FA_253: FA port map(pp(80), pp(57), pp(34), sum(252), carry(252));
	FA_254: FA port map(pp(11), carry(134), carry(133), sum(253), carry(253));
	FA_255: FA port map(sum(135), sum(136), sum(137), sum(254), carry(254));
	FA_256: FA port map(pp(35), pp(12), carry(137), sum(255), carry(255));
	FA_257: FA port map(carry(136), carry(135), sum(138), sum(256), carry(256));
	FA_258: FA port map(sum(139), sum(140), sum(141), sum(257), carry(257));
	FA_259: FA port map(sum(30), carry(141), carry(140), sum(258), carry(258));
	FA_260: FA port map(carry(139), carry(138), sum(142), sum(259), carry(259));
	FA_261: FA port map(sum(143), sum(144), sum(145), sum(260), carry(260));
	FA_262: FA port map(sum(32), carry(145), carry(144), sum(261), carry(261));
	FA_263: FA port map(carry(143), carry(142), sum(146), sum(262), carry(262));
	FA_264: FA port map(sum(147), sum(148), sum(149), sum(263), carry(263));
	FA_265: FA port map(sum(35), carry(149), carry(148), sum(264), carry(264));
	FA_266: FA port map(carry(147), carry(146), sum(150), sum(265), carry(265));
	FA_267: FA port map(sum(151), sum(152), sum(153), sum(266), carry(266));
	FA_268: FA port map(sum(39), carry(153), carry(152), sum(267), carry(267));
	FA_269: FA port map(carry(151), carry(150), sum(154), sum(268), carry(268));
	FA_270: FA port map(sum(155), sum(156), sum(157), sum(269), carry(269));
	FA_271: FA port map(sum(44), carry(157), carry(156), sum(270), carry(270));
	FA_272: FA port map(carry(155), carry(154), sum(158), sum(271), carry(271));
	FA_273: FA port map(sum(159), sum(160), sum(161), sum(272), carry(272));
	FA_274: FA port map(sum(50), carry(161), carry(160), sum(273), carry(273));
	FA_275: FA port map(carry(159), carry(158), sum(162), sum(274), carry(274));
	FA_276: FA port map(sum(163), sum(164), sum(165), sum(275), carry(275));
	FA_277: FA port map(sum(56), carry(165), carry(164), sum(276), carry(276));
	FA_278: FA port map(carry(163), carry(162), sum(166), sum(277), carry(277));
	FA_279: FA port map(sum(167), sum(168), sum(169), sum(278), carry(278));
	FA_280: FA port map(sum(62), carry(169), carry(168), sum(279), carry(279));
	FA_281: FA port map(carry(167), carry(166), sum(170), sum(280), carry(280));
	FA_282: FA port map(sum(171), sum(172), sum(173), sum(281), carry(281));
	FA_283: FA port map(sum(68), carry(173), carry(172), sum(282), carry(282));
	FA_284: FA port map(carry(171), carry(170), sum(174), sum(283), carry(283));
	FA_285: FA port map(sum(175), sum(176), sum(177), sum(284), carry(284));
	FA_286: FA port map(sum(74), carry(177), carry(176), sum(285), carry(285));
	FA_287: FA port map(carry(175), carry(174), sum(178), sum(286), carry(286));
	FA_288: FA port map(sum(179), sum(180), sum(181), sum(287), carry(287));
	FA_289: FA port map(sum(80), carry(181), carry(180), sum(288), carry(288));
	FA_290: FA port map(carry(179), carry(178), sum(182), sum(289), carry(289));
	FA_291: FA port map(sum(183), sum(184), sum(185), sum(290), carry(290));
	FA_292: FA port map(sum(86), carry(185), carry(184), sum(291), carry(291));
	FA_293: FA port map(carry(183), carry(182), sum(186), sum(292), carry(292));
	FA_294: FA port map(sum(187), sum(188), sum(189), sum(293), carry(293));
	FA_295: FA port map(sum(92), carry(189), carry(188), sum(294), carry(294));
	FA_296: FA port map(carry(187), carry(186), sum(190), sum(295), carry(295));
	FA_297: FA port map(sum(191), sum(192), sum(193), sum(296), carry(296));
	FA_298: FA port map(sum(98), carry(193), carry(192), sum(297), carry(297));
	FA_299: FA port map(carry(191), carry(190), sum(194), sum(298), carry(298));
	FA_300: FA port map(sum(195), sum(196), sum(197), sum(299), carry(299));
	FA_301: FA port map(sum(104), carry(197), carry(196), sum(300), carry(300));
	FA_302: FA port map(carry(195), carry(194), sum(198), sum(301), carry(301));
	FA_303: FA port map(sum(199), sum(200), sum(201), sum(302), carry(302));
	FA_304: FA port map(sum(110), carry(201), carry(200), sum(303), carry(303));
	FA_305: FA port map(carry(199), carry(198), sum(202), sum(304), carry(304));
	FA_306: FA port map(sum(203), sum(204), sum(205), sum(305), carry(305));
	FA_307: FA port map(sum(116), carry(205), carry(204), sum(306), carry(306));
	FA_308: FA port map(carry(203), carry(202), sum(206), sum(307), carry(307));
	FA_309: FA port map(sum(207), sum(208), sum(209), sum(308), carry(308));
	FA_310: FA port map(sum(121), carry(209), carry(208), sum(309), carry(309));
	FA_311: FA port map(carry(207), carry(206), sum(210), sum(310), carry(310));
	FA_312: FA port map(sum(211), sum(212), sum(213), sum(311), carry(311));
	FA_313: FA port map(sum(125), carry(213), carry(212), sum(312), carry(312));
	FA_314: FA port map(carry(211), carry(210), sum(214), sum(313), carry(313));
	FA_315: FA port map(sum(215), sum(216), sum(217), sum(314), carry(314));
	FA_316: FA port map(sum(128), carry(217), carry(216), sum(315), carry(315));
	FA_317: FA port map(carry(215), carry(214), sum(218), sum(316), carry(316));
	FA_318: FA port map(sum(219), sum(220), sum(221), sum(317), carry(317));
	FA_319: FA port map(sum(130), carry(221), carry(220), sum(318), carry(318));
	FA_320: FA port map(carry(219), carry(218), sum(222), sum(319), carry(319));
	FA_321: FA port map(sum(223), sum(224), sum(225), sum(320), carry(320));
	FA_322: FA port map(sum(131), carry(225), carry(224), sum(321), carry(321));
	FA_323: FA port map(carry(223), carry(222), sum(226), sum(322), carry(322));
	FA_324: FA port map(sum(227), sum(228), sum(229), sum(323), carry(323));
	FA_325: FA port map(carry(131), carry(229), carry(228), sum(324), carry(324));
	FA_326: FA port map(carry(227), carry(226), sum(230), sum(325), carry(325));
	FA_327: FA port map(sum(231), sum(232), sum(233), sum(326), carry(326));
	FA_328: FA port map(pp(358), pp(335), carry(233), sum(327), carry(327));
	FA_329: FA port map(carry(232), carry(231), carry(230), sum(328), carry(328));
	FA_330: FA port map(sum(234), sum(235), sum(236), sum(329), carry(329));
	FA_331: FA port map(pp(428), pp(405), pp(382), sum(330), carry(330));
	FA_332: FA port map(pp(359), carry(236), carry(235), sum(331), carry(331));
	FA_333: FA port map(carry(234), sum(237), sum(238), sum(332), carry(332));
	FA_334: FA port map(pp(498), pp(475), pp(452), sum(333), carry(333));
	FA_335: FA port map(pp(429), pp(406), pp(383), sum(334), carry(334));
	FA_336: FA port map(carry(238), carry(237), sum(239), sum(335), carry(335));
	FA_337: FA port map(pp(568), pp(545), pp(522), sum(336), carry(336));
	FA_338: FA port map(pp(499), pp(476), pp(453), sum(337), carry(337));
	FA_339: FA port map(pp(430), pp(407), carry(239), sum(338), carry(338));
	FA_340: FA port map(pp(569), pp(546), pp(523), sum(339), carry(339));
	FA_341: FA port map(pp(500), pp(477), pp(454), sum(340), carry(340));
	FA_342: FA port map(pp(570), pp(547), pp(524), sum(341), carry(341));
	
	-- Stage J = 3; d_3 = 4
	-- HAs ALLOCATED: 2 (21 TOTAL)
	-- FAs ALLOCATED: 76 (399 TOTAL)
	HA_343: HA port map(pp(96), pp(73), sum(342), carry(342));
	FA_344: FA port map(pp(120), pp(97), pp(74), sum(343), carry(343));
	HA_345: HA port map(pp(51), pp(28), sum(344), carry(344));
	FA_346: FA port map(pp(98), pp(75), pp(52), sum(345), carry(345));
	FA_347: FA port map(pp(29), pp(6), sum(240), sum(346), carry(346));
	FA_348: FA port map(pp(53), pp(30), pp(7), sum(347), carry(347));
	FA_349: FA port map(carry(240), sum(241), sum(242), sum(348), carry(348));
	FA_350: FA port map(pp(8), carry(242), carry(241), sum(349), carry(349));
	FA_351: FA port map(sum(243), sum(244), sum(245), sum(350), carry(350));
	FA_352: FA port map(carry(245), carry(244), carry(243), sum(351), carry(351));
	FA_353: FA port map(sum(246), sum(247), sum(248), sum(352), carry(352));
	FA_354: FA port map(carry(248), carry(247), carry(246), sum(353), carry(353));
	FA_355: FA port map(sum(249), sum(250), sum(251), sum(354), carry(354));
	FA_356: FA port map(carry(251), carry(250), carry(249), sum(355), carry(355));
	FA_357: FA port map(sum(252), sum(253), sum(254), sum(356), carry(356));
	FA_358: FA port map(carry(254), carry(253), carry(252), sum(357), carry(357));
	FA_359: FA port map(sum(255), sum(256), sum(257), sum(358), carry(358));
	FA_360: FA port map(carry(257), carry(256), carry(255), sum(359), carry(359));
	FA_361: FA port map(sum(258), sum(259), sum(260), sum(360), carry(360));
	FA_362: FA port map(carry(260), carry(259), carry(258), sum(361), carry(361));
	FA_363: FA port map(sum(261), sum(262), sum(263), sum(362), carry(362));
	FA_364: FA port map(carry(263), carry(262), carry(261), sum(363), carry(363));
	FA_365: FA port map(sum(264), sum(265), sum(266), sum(364), carry(364));
	FA_366: FA port map(carry(266), carry(265), carry(264), sum(365), carry(365));
	FA_367: FA port map(sum(267), sum(268), sum(269), sum(366), carry(366));
	FA_368: FA port map(carry(269), carry(268), carry(267), sum(367), carry(367));
	FA_369: FA port map(sum(270), sum(271), sum(272), sum(368), carry(368));
	FA_370: FA port map(carry(272), carry(271), carry(270), sum(369), carry(369));
	FA_371: FA port map(sum(273), sum(274), sum(275), sum(370), carry(370));
	FA_372: FA port map(carry(275), carry(274), carry(273), sum(371), carry(371));
	FA_373: FA port map(sum(276), sum(277), sum(278), sum(372), carry(372));
	FA_374: FA port map(carry(278), carry(277), carry(276), sum(373), carry(373));
	FA_375: FA port map(sum(279), sum(280), sum(281), sum(374), carry(374));
	FA_376: FA port map(carry(281), carry(280), carry(279), sum(375), carry(375));
	FA_377: FA port map(sum(282), sum(283), sum(284), sum(376), carry(376));
	FA_378: FA port map(carry(284), carry(283), carry(282), sum(377), carry(377));
	FA_379: FA port map(sum(285), sum(286), sum(287), sum(378), carry(378));
	FA_380: FA port map(carry(287), carry(286), carry(285), sum(379), carry(379));
	FA_381: FA port map(sum(288), sum(289), sum(290), sum(380), carry(380));
	FA_382: FA port map(carry(290), carry(289), carry(288), sum(381), carry(381));
	FA_383: FA port map(sum(291), sum(292), sum(293), sum(382), carry(382));
	FA_384: FA port map(carry(293), carry(292), carry(291), sum(383), carry(383));
	FA_385: FA port map(sum(294), sum(295), sum(296), sum(384), carry(384));
	FA_386: FA port map(carry(296), carry(295), carry(294), sum(385), carry(385));
	FA_387: FA port map(sum(297), sum(298), sum(299), sum(386), carry(386));
	FA_388: FA port map(carry(299), carry(298), carry(297), sum(387), carry(387));
	FA_389: FA port map(sum(300), sum(301), sum(302), sum(388), carry(388));
	FA_390: FA port map(carry(302), carry(301), carry(300), sum(389), carry(389));
	FA_391: FA port map(sum(303), sum(304), sum(305), sum(390), carry(390));
	FA_392: FA port map(carry(305), carry(304), carry(303), sum(391), carry(391));
	FA_393: FA port map(sum(306), sum(307), sum(308), sum(392), carry(392));
	FA_394: FA port map(carry(308), carry(307), carry(306), sum(393), carry(393));
	FA_395: FA port map(sum(309), sum(310), sum(311), sum(394), carry(394));
	FA_396: FA port map(carry(311), carry(310), carry(309), sum(395), carry(395));
	FA_397: FA port map(sum(312), sum(313), sum(314), sum(396), carry(396));
	FA_398: FA port map(carry(314), carry(313), carry(312), sum(397), carry(397));
	FA_399: FA port map(sum(315), sum(316), sum(317), sum(398), carry(398));
	FA_400: FA port map(carry(317), carry(316), carry(315), sum(399), carry(399));
	FA_401: FA port map(sum(318), sum(319), sum(320), sum(400), carry(400));
	FA_402: FA port map(carry(320), carry(319), carry(318), sum(401), carry(401));
	FA_403: FA port map(sum(321), sum(322), sum(323), sum(402), carry(402));
	FA_404: FA port map(carry(323), carry(322), carry(321), sum(403), carry(403));
	FA_405: FA port map(sum(324), sum(325), sum(326), sum(404), carry(404));
	FA_406: FA port map(carry(326), carry(325), carry(324), sum(405), carry(405));
	FA_407: FA port map(sum(327), sum(328), sum(329), sum(406), carry(406));
	FA_408: FA port map(carry(329), carry(328), carry(327), sum(407), carry(407));
	FA_409: FA port map(sum(330), sum(331), sum(332), sum(408), carry(408));
	FA_410: FA port map(carry(332), carry(331), carry(330), sum(409), carry(409));
	FA_411: FA port map(sum(333), sum(334), sum(335), sum(410), carry(410));
	FA_412: FA port map(carry(335), carry(334), carry(333), sum(411), carry(411));
	FA_413: FA port map(sum(336), sum(337), sum(338), sum(412), carry(412));
	FA_414: FA port map(pp(431), carry(338), carry(337), sum(413), carry(413));
	FA_415: FA port map(carry(336), sum(339), sum(340), sum(414), carry(414));
	FA_416: FA port map(pp(501), pp(478), pp(455), sum(415), carry(415));
	FA_417: FA port map(carry(340), carry(339), sum(341), sum(416), carry(416));
	FA_418: FA port map(pp(571), pp(548), pp(525), sum(417), carry(417));
	FA_419: FA port map(pp(502), pp(479), carry(341), sum(418), carry(418));
	FA_420: FA port map(pp(572), pp(549), pp(526), sum(419), carry(419));
	
	-- Stage J = 2; d_2 = 3
	-- HAs ALLOCATED: 1 (22 TOTAL)
	-- FAs ALLOCATED: 41 (440 TOTAL)
	HA_421: HA port map(pp(72), pp(49), sum(420), carry(420));
	FA_422: FA port map(pp(50), pp(27), pp(4), sum(421), carry(421));
	FA_423: FA port map(pp(5), carry(342), sum(343), sum(422), carry(422));
	FA_424: FA port map(carry(344), carry(343), sum(345), sum(423), carry(423));
	FA_425: FA port map(carry(346), carry(345), sum(347), sum(424), carry(424));
	FA_426: FA port map(carry(348), carry(347), sum(349), sum(425), carry(425));
	FA_427: FA port map(carry(350), carry(349), sum(351), sum(426), carry(426));
	FA_428: FA port map(carry(352), carry(351), sum(353), sum(427), carry(427));
	FA_429: FA port map(carry(354), carry(353), sum(355), sum(428), carry(428));
	FA_430: FA port map(carry(356), carry(355), sum(357), sum(429), carry(429));
	FA_431: FA port map(carry(358), carry(357), sum(359), sum(430), carry(430));
	FA_432: FA port map(carry(360), carry(359), sum(361), sum(431), carry(431));
	FA_433: FA port map(carry(362), carry(361), sum(363), sum(432), carry(432));
	FA_434: FA port map(carry(364), carry(363), sum(365), sum(433), carry(433));
	FA_435: FA port map(carry(366), carry(365), sum(367), sum(434), carry(434));
	FA_436: FA port map(carry(368), carry(367), sum(369), sum(435), carry(435));
	FA_437: FA port map(carry(370), carry(369), sum(371), sum(436), carry(436));
	FA_438: FA port map(carry(372), carry(371), sum(373), sum(437), carry(437));
	FA_439: FA port map(carry(374), carry(373), sum(375), sum(438), carry(438));
	FA_440: FA port map(carry(376), carry(375), sum(377), sum(439), carry(439));
	FA_441: FA port map(carry(378), carry(377), sum(379), sum(440), carry(440));
	FA_442: FA port map(carry(380), carry(379), sum(381), sum(441), carry(441));
	FA_443: FA port map(carry(382), carry(381), sum(383), sum(442), carry(442));
	FA_444: FA port map(carry(384), carry(383), sum(385), sum(443), carry(443));
	FA_445: FA port map(carry(386), carry(385), sum(387), sum(444), carry(444));
	FA_446: FA port map(carry(388), carry(387), sum(389), sum(445), carry(445));
	FA_447: FA port map(carry(390), carry(389), sum(391), sum(446), carry(446));
	FA_448: FA port map(carry(392), carry(391), sum(393), sum(447), carry(447));
	FA_449: FA port map(carry(394), carry(393), sum(395), sum(448), carry(448));
	FA_450: FA port map(carry(396), carry(395), sum(397), sum(449), carry(449));
	FA_451: FA port map(carry(398), carry(397), sum(399), sum(450), carry(450));
	FA_452: FA port map(carry(400), carry(399), sum(401), sum(451), carry(451));
	FA_453: FA port map(carry(402), carry(401), sum(403), sum(452), carry(452));
	FA_454: FA port map(carry(404), carry(403), sum(405), sum(453), carry(453));
	FA_455: FA port map(carry(406), carry(405), sum(407), sum(454), carry(454));
	FA_456: FA port map(carry(408), carry(407), sum(409), sum(455), carry(455));
	FA_457: FA port map(carry(410), carry(409), sum(411), sum(456), carry(456));
	FA_458: FA port map(carry(412), carry(411), sum(413), sum(457), carry(457));
	FA_459: FA port map(carry(414), carry(413), sum(415), sum(458), carry(458));
	FA_460: FA port map(carry(416), carry(415), sum(417), sum(459), carry(459));
	FA_461: FA port map(pp(503), carry(418), carry(417), sum(460), carry(460));
	FA_462: FA port map(pp(573), pp(550), pp(527), sum(461), carry(461));
	
	-- Stage J = 1; d_1 = 2
	-- HAs ALLOCATED: 1 (23 TOTAL)
	-- FAs ALLOCATED: 43 (483 TOTAL)
	HA_463: HA port map(pp(48), pp(25), sum(462), carry(462));
	FA_464: FA port map(pp(26), pp(3), sum(420), sum(463), carry(463));
	FA_465: FA port map(sum(342), carry(420), sum(421), sum(464), carry(464));
	FA_466: FA port map(sum(344), carry(421), sum(422), sum(465), carry(465));
	FA_467: FA port map(sum(346), carry(422), sum(423), sum(466), carry(466));
	FA_468: FA port map(sum(348), carry(423), sum(424), sum(467), carry(467));
	FA_469: FA port map(sum(350), carry(424), sum(425), sum(468), carry(468));
	FA_470: FA port map(sum(352), carry(425), sum(426), sum(469), carry(469));
	FA_471: FA port map(sum(354), carry(426), sum(427), sum(470), carry(470));
	FA_472: FA port map(sum(356), carry(427), sum(428), sum(471), carry(471));
	FA_473: FA port map(sum(358), carry(428), sum(429), sum(472), carry(472));
	FA_474: FA port map(sum(360), carry(429), sum(430), sum(473), carry(473));
	FA_475: FA port map(sum(362), carry(430), sum(431), sum(474), carry(474));
	FA_476: FA port map(sum(364), carry(431), sum(432), sum(475), carry(475));
	FA_477: FA port map(sum(366), carry(432), sum(433), sum(476), carry(476));
	FA_478: FA port map(sum(368), carry(433), sum(434), sum(477), carry(477));
	FA_479: FA port map(sum(370), carry(434), sum(435), sum(478), carry(478));
	FA_480: FA port map(sum(372), carry(435), sum(436), sum(479), carry(479));
	FA_481: FA port map(sum(374), carry(436), sum(437), sum(480), carry(480));
	FA_482: FA port map(sum(376), carry(437), sum(438), sum(481), carry(481));
	FA_483: FA port map(sum(378), carry(438), sum(439), sum(482), carry(482));
	FA_484: FA port map(sum(380), carry(439), sum(440), sum(483), carry(483));
	FA_485: FA port map(sum(382), carry(440), sum(441), sum(484), carry(484));
	FA_486: FA port map(sum(384), carry(441), sum(442), sum(485), carry(485));
	FA_487: FA port map(sum(386), carry(442), sum(443), sum(486), carry(486));
	FA_488: FA port map(sum(388), carry(443), sum(444), sum(487), carry(487));
	FA_489: FA port map(sum(390), carry(444), sum(445), sum(488), carry(488));
	FA_490: FA port map(sum(392), carry(445), sum(446), sum(489), carry(489));
	FA_491: FA port map(sum(394), carry(446), sum(447), sum(490), carry(490));
	FA_492: FA port map(sum(396), carry(447), sum(448), sum(491), carry(491));
	FA_493: FA port map(sum(398), carry(448), sum(449), sum(492), carry(492));
	FA_494: FA port map(sum(400), carry(449), sum(450), sum(493), carry(493));
	FA_495: FA port map(sum(402), carry(450), sum(451), sum(494), carry(494));
	FA_496: FA port map(sum(404), carry(451), sum(452), sum(495), carry(495));
	FA_497: FA port map(sum(406), carry(452), sum(453), sum(496), carry(496));
	FA_498: FA port map(sum(408), carry(453), sum(454), sum(497), carry(497));
	FA_499: FA port map(sum(410), carry(454), sum(455), sum(498), carry(498));
	FA_500: FA port map(sum(412), carry(455), sum(456), sum(499), carry(499));
	FA_501: FA port map(sum(414), carry(456), sum(457), sum(500), carry(500));
	FA_502: FA port map(sum(416), carry(457), sum(458), sum(501), carry(501));
	FA_503: FA port map(sum(418), carry(458), sum(459), sum(502), carry(502));
	FA_504: FA port map(sum(419), carry(459), sum(460), sum(503), carry(503));
	FA_505: FA port map(carry(419), carry(460), sum(461), sum(504), carry(504));
	FA_506: FA port map(pp(574), pp(551), carry(461), sum(505), carry(505));
	

	-- FINAL ADDER
	PROD(0) <= pp(0);
	final_adder_op1(45 downto 0) <= pp(575) & carry(504) & carry(503) & carry(502) & carry(501) & carry(500) & carry(499) & carry(498) & carry(497) & carry(496) & carry(495) & carry(494) & carry(493) & carry(492) & carry(491) & carry(490) & carry(489) & carry(488) & carry(487) & carry(486) & carry(485) & carry(484) & carry(483) & carry(482) & carry(481) & carry(480) & carry(479) & carry(478) & carry(477) & carry(476) & carry(475) & carry(474) & carry(473) & carry(472) & carry(471) & carry(470) & carry(469) & carry(468) & carry(467) & carry(466) & carry(465) & carry(464) & carry(463) & carry(462) & pp(2) & pp(24);
	final_adder_op2(45 downto 0) <= carry(505) & sum(505) & sum(504) & sum(503) & sum(502) & sum(501) & sum(500) & sum(499) & sum(498) & sum(497) & sum(496) & sum(495) & sum(494) & sum(493) & sum(492) & sum(491) & sum(490) & sum(489) & sum(488) & sum(487) & sum(486) & sum(485) & sum(484) & sum(483) & sum(482) & sum(481) & sum(480) & sum(479) & sum(478) & sum(477) & sum(476) & sum(475) & sum(474) & sum(473) & sum(472) & sum(471) & sum(470) & sum(469) & sum(468) & sum(467) & sum(466) & sum(465) & sum(464) & sum(463) & sum(462) & pp(1);
	final_adder_op1(46) <= '0';
	final_adder_op2(46) <= '0';
	final_adder_sum <= to_integer(unsigned(final_adder_op1)) + to_integer(unsigned(final_adder_op2));
	PROD(47 downto 1) <= std_logic_vector(to_unsigned(final_adder_sum,47));

end architecture;