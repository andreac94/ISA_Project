package integer_array is
    type int_array is array(integer range <>) of integer;
end package integer_array;
